// Execute test bench module
module execute_tb ();

  // Parameters
  parameter CNT_TESTS = 100;  // cnt of tests

  // Test bench variables
  logic clk, reset_tb;
  logic [63 : 0] PCBranch_E_expected, aluResult_E_expected, writeData_E_expected;
  logic zero_E_expected;

  int test_number, cnt_errors;
  logic [453 : 0] test[0 : CNT_TESTS-1];
  // {{AluSrc}, {AluControl}, {PC_E}, {signImm_E}, {readData1_E}, {readData2_E}, {PCBranch_E_expected}, {aluResult_E_expected}, {writeData_E_expected}, {zero_E_expected}}

  // Module connections
  logic AluSrc, zero_E;
  logic [3 : 0] AluControl;
  logic [63 : 0] PC_E, signImm_E, readData1_E, readData2_E, PCBranch_E, aluResult_E, writeData_E;

  execute dut (
      .AluSrc(AluSrc),
      .AluControl(AluControl),
      .PC_E(PC_E),
      .signImm_E(signImm_E),
      .readData1_E(readData1_E),
      .readData2_E(readData2_E),
      .PCBranch_E(PCBranch_E),
      .aluResult_E(aluResult_E),
      .writeData_E(writeData_E),
      .zero_E(zero_E)
  );

  // Clock generation with 10ns period
  always begin
    clk = 1;
    #5ns;
    clk = 0;
    #5ns;
  end

  initial begin
    // Init tests
    test_number = 0;
    cnt_errors = 0;

    test = {
      {
        {1'd1},
        {4'd1},
        {64'd275899981746774790},
        {64'd1146357998626863111},
        {64'd417007973947494494},
        {64'd290168482088084069},
        {64'd4861331976254227234},
        {64'd1146639509341206623},
        {64'd290168482088084069},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd560809363472268348},
        {64'd1086815724955799638},
        {64'd791603134059380040},
        {64'd443955406591393154},
        {64'd4908072263295466900},
        {64'd1152209021055139166},
        {64'd443955406591393154},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd780331085967984627},
        {64'd508225762828702171},
        {64'd1127686399091378860},
        {64'd1079334227989712615},
        {64'd2813234137282793311},
        {64'd505547209291399304},
        {64'd1079334227989712615},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd695426852230382782},
        {64'd393282134813786452},
        {64'd532276753602227935},
        {64'd261213995781211471},
        {64'd2268555391485528590},
        {64'd537967845418332127},
        {64'd261213995781211471},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd736093754794182240},
        {64'd1003195744507934607},
        {64'd974456296342379981},
        {64'd1115026736238234457},
        {64'd4748876732825920668},
        {64'd1115026736238234457},
        {64'd1115026736238234457},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd627544731619043598},
        {64'd385128650287974267},
        {64'd91523881260785684},
        {64'd123940227453340073},
        {64'd2168059332770940666},
        {64'd386580040634050431},
        {64'd123940227453340073},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd630044586087911607},
        {64'd690212882881701560},
        {64'd3100836379041554},
        {64'd490174023508158029},
        {64'd3390896117614717847},
        {64'd690212882881701560},
        {64'd490174023508158029},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd535040534797432328},
        {64'd572613525127545460},
        {64'd507846478024118271},
        {64'd713121694943710190},
        {64'd2825494635307614168},
        {64'd504421463853335156},
        {64'd713121694943710190},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd793948544465316899},
        {64'd19350433455582208},
        {64'd273513854920686606},
        {64'd335908015352833116},
        {64'd871350278287645731},
        {64'd292864288376268814},
        {64'd335908015352833116},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd14616297492838228},
        {64'd1134982342437728350},
        {64'd98388997430521492},
        {64'd1050619260381204426},
        {64'd4554545667243751628},
        {64'd1050619260381204426},
        {64'd1050619260381204426},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd350604512921165627},
        {64'd703018173509345534},
        {64'd300638415632515183},
        {64'd607224119094326764},
        {64'd3162677206958547763},
        {64'd23131897462894},
        {64'd607224119094326764},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd648022744817110269},
        {64'd588010465796643684},
        {64'd67422489384660151},
        {64'd491761106988897620},
        {64'd3000064608003685005},
        {64'd491761106988897620},
        {64'd491761106988897620},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd822593250848530524},
        {64'd878608095165024603},
        {64'd331620452017095461},
        {64'd28780789398848009},
        {64'd4337025631508628936},
        {64'd302839662618247452},
        {64'd28780789398848009},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd738416654991249802},
        {64'd550647299411546728},
        {64'd283613051013701000},
        {64'd992270869193736727},
        {64'd2941005852637436714},
        {64'd571916321360846824},
        {64'd992270869193736727},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd567363897597520658},
        {64'd131720619578627738},
        {64'd829175074006215547},
        {64'd456531573305056694},
        {64'd1094246375912031610},
        {64'd372643500701158853},
        {64'd456531573305056694},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd84963837130065931},
        {64'd349698210751673725},
        {64'd1024413202427644553},
        {64'd1021185305924167092},
        {64'd1483756680136760831},
        {64'd293402621797007369},
        {64'd1021185305924167092},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd449588735098673247},
        {64'd265727246895323808},
        {64'd496737682936494336},
        {64'd1095737244521803015},
        {64'd1512497722679968479},
        {64'd1592474927458297351},
        {64'd1095737244521803015},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd825221091594656384},
        {64'd1095741053695843895},
        {64'd692837975977287035},
        {64'd492085617346702144},
        {64'd5208185306378031964},
        {64'd1184923593323989179},
        {64'd492085617346702144},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd48606430248752046},
        {64'd90539929078548686},
        {64'd570385732746553284},
        {64'd119678457820111415},
        {64'd410766146562946790},
        {64'd570671743554775031},
        {64'd119678457820111415},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd683353024891835270},
        {64'd1053226656510633735},
        {64'd10874906354945493},
        {64'd587296358288181977},
        {64'd4896259650934370210},
        {64'd1062834924123975639},
        {64'd587296358288181977},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd502434407369840338},
        {64'd654829103297569279},
        {64'd156495987410662235},
        {64'd790878865902613692},
        {64'd3121750820560117454},
        {64'd790878865902613692},
        {64'd790878865902613692},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd1012070287809094604},
        {64'd483341090482292628},
        {64'd1142807559916959076},
        {64'd713943308184603321},
        {64'd2945434649738265116},
        {64'd1152144612668684276},
        {64'd713943308184603321},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd832231367132619876},
        {64'd997206744208682347},
        {64'd446550633026245295},
        {64'd444139702044595752},
        {64'd4821058343967349264},
        {64'd1150387608655757295},
        {64'd444139702044595752},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd337132479512866020},
        {64'd363562185325618564},
        {64'd101593663745081811},
        {64'd221058537083930738},
        {64'd1791381220815340276},
        {64'd18327279200370702689},
        {64'd221058537083930738},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd53997849180224586},
        {64'd1023962611639106403},
        {64'd838308817520562486},
        {64'd1075915243241177868},
        {64'd4149848295736650198},
        {64'd729653515089350946},
        {64'd1075915243241177868},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd927777055475948315},
        {64'd1073689159693010433},
        {64'd637758216571836713},
        {64'd207072713736922155},
        {64'd5222533694247990047},
        {64'd1080802038074957609},
        {64'd207072713736922155},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd427981837430653748},
        {64'd63785584533024260},
        {64'd898251533437188842},
        {64'd317157228970134246},
        {64'd683124175562750788},
        {64'd581094304467054596},
        {64'd317157228970134246},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd746425135871551828},
        {64'd903289679994987195},
        {64'd280858537801578080},
        {64'd245967566702009487},
        {64'd4359583855851500608},
        {64'd243698033538651136},
        {64'd245967566702009487},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd240315894690958431},
        {64'd1002607669530085280},
        {64'd1055638316964331030},
        {64'd143206706099814954},
        {64'd4250746572811299551},
        {64'd909833038712538624},
        {64'd143206706099814954},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd361519145694254601},
        {64'd112570993416474595},
        {64'd1054445822201868808},
        {64'd11431499853174359},
        {64'd811803119360152981},
        {64'd1043014322348694449},
        {64'd11431499853174359},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd345873591510464484},
        {64'd172150533461421328},
        {64'd1022103174697045994},
        {64'd408399014252971974},
        {64'd1034475725356149796},
        {64'd408399014252971974},
        {64'd408399014252971974},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd870530475273287314},
        {64'd180201444928259912},
        {64'd1017946893915769981},
        {64'd423863973786591753},
        {64'd1591336254986326962},
        {64'd594082920129178228},
        {64'd423863973786591753},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd183806536705535283},
        {64'd943503058793357598},
        {64'd535762376489349798},
        {64'd454666611194828844},
        {64'd3957818771878965675},
        {64'd1479265435282707396},
        {64'd454666611194828844},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd489452135262500359},
        {64'd720942297253462869},
        {64'd162013147177498229},
        {64'd996549582525998037},
        {64'd3373221324276351835},
        {64'd17612207638361051808},
        {64'd996549582525998037},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd206297714561374278},
        {64'd55684996594435655},
        {64'd975130522794990646},
        {64'd790063936243571646},
        {64'd429037700939116898},
        {64'd612590714131585078},
        {64'd790063936243571646},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd758031223640297279},
        {64'd712022199616142026},
        {64'd773371864695859393},
        {64'd490541505774200565},
        {64'd3606120022104865383},
        {64'd183100039323721921},
        {64'd490541505774200565},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd172597629290264975},
        {64'd133366409688245907},
        {64'd205498203234650698},
        {64'd1011464410819244655},
        {64'd706063268043248603},
        {64'd1070576364079086191},
        {64'd1011464410819244655},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd396591846936414043},
        {64'd550946586539517485},
        {64'd1015998066520835315},
        {64'd61516834974626498},
        {64'd2600378193094483983},
        {64'd1077514901495461813},
        {64'd61516834974626498},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd8988875185501022},
        {64'd960320253047926838},
        {64'd332844953834408476},
        {64'd323642033338484037},
        {64'd3850269887377208374},
        {64'd323642033338484037},
        {64'd323642033338484037},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd821978214028015560},
        {64'd386076487913717228},
        {64'd264504401106844627},
        {64'd506541609155016786},
        {64'd2366284165682884472},
        {64'd650580889020561855},
        {64'd506541609155016786},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd698296927504805769},
        {64'd511872762092337269},
        {64'd582611692593249655},
        {64'd275211241139853529},
        {64'd2745787975874154845},
        {64'd511872762092337269},
        {64'd275211241139853529},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd609923247257659993},
        {64'd825311591562875548},
        {64'd808717145004402798},
        {64'd757650117468179018},
        {64'd3911169613509162185},
        {64'd720895640623728714},
        {64'd757650117468179018},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd344871138391749298},
        {64'd490951676866572007},
        {64'd847518908774563063},
        {64'd5745545478741951},
        {64'd2308677845858037326},
        {64'd853264454253305014},
        {64'd5745545478741951},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd204363087088465424},
        {64'd885502219514464382},
        {64'd673893907951618590},
        {64'd75257900925178434},
        {64'd3746371965146322952},
        {64'd885502219514464382},
        {64'd75257900925178434},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd656449600917015319},
        {64'd12367672783375992},
        {64'd742706636700583454},
        {64'd27834663323888226},
        {64'd705920292050519287},
        {64'd18721659378467330},
        {64'd27834663323888226},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd422438424199615195},
        {64'd35146518124988234},
        {64'd574702688505073864},
        {64'd524923384850614228},
        {64'd563024496699568131},
        {64'd33989204288372808},
        {64'd524923384850614228},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd709423558383267009},
        {64'd368598260640470822},
        {64'd390083498529457747},
        {64'd301238821602833757},
        {64'd2183816600945150297},
        {64'd758681759169928569},
        {64'd301238821602833757},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd100535760635044553},
        {64'd1072494180515896870},
        {64'd936734734941474267},
        {64'd890180050701997266},
        {64'd4390512482698632033},
        {64'd890180050701997266},
        {64'd890180050701997266},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd588250433312659257},
        {64'd835893782013346528},
        {64'd208132357251399581},
        {64'd668484539117230090},
        {64'd3931825561366045369},
        {64'd18699413583583240},
        {64'd668484539117230090},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd415981874735463247},
        {64'd1117398165730229022},
        {64'd460273888819429716},
        {64'd432719396642341616},
        {64'd4885574537656379335},
        {64'd1117398165730229022},
        {64'd432719396642341616},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd761029197438090041},
        {64'd675948536176010095},
        {64'd1045413879164782250},
        {64'd448108388471274559},
        {64'd3464823342142130421},
        {64'd1061176565925412543},
        {64'd448108388471274559},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd61847399355904863},
        {64'd52045841408882466},
        {64'd793823570080884828},
        {64'd177711561669138070},
        {64'd270030764991434727},
        {64'd52045841408882466},
        {64'd177711561669138070},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd505899392868168167},
        {64'd835463528513442992},
        {64'd536308259789832},
        {64'd324993867164287914},
        {64'd3847753506921940135},
        {64'd17611816853455898456},
        {64'd324993867164287914},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd438106545851581041},
        {64'd926349670186608949},
        {64'd318018729312047562},
        {64'd806965183182834296},
        {64'd4143505226598016837},
        {64'd9218344151449672},
        {64'd806965183182834296},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd1137694605370527370},
        {64'd256216958325719716},
        {64'd1048268509137460719},
        {64'd139795144961797855},
        {64'd2162562438673406234},
        {64'd908473364175662864},
        {64'd139795144961797855},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd481548084006461633},
        {64'd1034272919533326623},
        {64'd82693311032202439},
        {64'd859086615722732435},
        {64'd4618639762139768125},
        {64'd1116966230565529062},
        {64'd859086615722732435},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd751663586319233082},
        {64'd661579426681436358},
        {64'd169644103021746177},
        {64'd395145790193991499},
        {64'd3397981293044978514},
        {64'd18221242386537306294},
        {64'd395145790193991499},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd917251240947251642},
        {64'd504139287522263264},
        {64'd45141007843249327},
        {64'd1054819756460082559},
        {64'd2933808391036304698},
        {64'd17437065325092718384},
        {64'd1054819756460082559},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd1120269218192893563},
        {64'd1115993475107334769},
        {64'd1152318057278243545},
        {64'd616759224756367941},
        {64'd5584243118622232639},
        {64'd535558832521875604},
        {64'd616759224756367941},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd249330614211506046},
        {64'd919986247500930588},
        {64'd80509137111123770},
        {64'd146105669535696297},
        {64'd3929275604215228398},
        {64'd18381147541284979089},
        {64'd146105669535696297},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd84293540099113048},
        {64'd594914848763814233},
        {64'd174383940095647469},
        {64'd212285389870819083},
        {64'd2463952935154369980},
        {64'd18408842623934380002},
        {64'd212285389870819083},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd542847240041253354},
        {64'd231556402973452764},
        {64'd643667746842831010},
        {64'd964181735564925074},
        {64'd1469072851935064410},
        {64'd412111343869378246},
        {64'd964181735564925074},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd1019117573072434683},
        {64'd967025618671512865},
        {64'd568309650173502551},
        {64'd1068880188955826075},
        {64'd4887220047758486143},
        {64'd18048028105211541302},
        {64'd1068880188955826075},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd1063136943314290658},
        {64'd439434016136489445},
        {64'd908111214681307076},
        {64'd1061878368459771965},
        {64'd2820873007860248438},
        {64'd1052556978874351589},
        {64'd1061878368459771965},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd980012907534982755},
        {64'd811155991557886503},
        {64'd993869562849057374},
        {64'd908466768123086783},
        {64'd4224636873766528767},
        {64'd1805025554406943877},
        {64'd908466768123086783},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd570797562185921377},
        {64'd626092778197131116},
        {64'd977915103139773429},
        {64'd802409504458842964},
        {64'd3075168674974445841},
        {64'd1780324607598616393},
        {64'd802409504458842964},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd173426364220889484},
        {64'd230446325298562220},
        {64'd415727974025023742},
        {64'd547676614405370648},
        {64'd1095211665415138364},
        {64'd573918647059698942},
        {64'd547676614405370648},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd443892723142259385},
        {64'd200753278763987907},
        {64'd703797939113269336},
        {64'd817426381263208544},
        {64'd1246905838198211013},
        {64'd200753278763987907},
        {64'd817426381263208544},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd257467357703654477},
        {64'd979478877765172990},
        {64'd420273695900906107},
        {64'd1049481051074920515},
        {64'd4175382868764346437},
        {64'd1140991768009847419},
        {64'd1049481051074920515},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd323025669870392558},
        {64'd343046629524241319},
        {64'd382639247113758616},
        {64'd700385339654795972},
        {64'd1695212187967357834},
        {64'd700385339654795972},
        {64'd700385339654795972},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd693785987289030215},
        {64'd17089116158488923},
        {64'd230616065066192091},
        {64'd514056137481131384},
        {64'd762142451922985907},
        {64'd18163304001294612323},
        {64'd514056137481131384},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd434889272584206343},
        {64'd643437248802293543},
        {64'd813782895745607374},
        {64'd178772254340677436},
        {64'd3008638267793380515},
        {64'd635010641404929938},
        {64'd178772254340677436},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd765333545470094875},
        {64'd396923319208219514},
        {64'd953762513943193044},
        {64'd461133886719099052},
        {64'd2353026822302972931},
        {64'd990360874700765182},
        {64'd461133886719099052},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd1123710680535973796},
        {64'd186652929411824845},
        {64'd750359269769968133},
        {64'd327141417034138385},
        {64'd1870322398183273176},
        {64'd144413986811557893},
        {64'd327141417034138385},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd766160755862033176},
        {64'd44744576839930889},
        {64'd341705775789146458},
        {64'd1046327969646802345},
        {64'd945139063221756732},
        {64'd44744576839930889},
        {64'd1046327969646802345},
        {1'd0}
      },
      {
        {1'd1},
        {4'd1},
        {64'd1080444516535496224},
        {64'd195834180266931850},
        {64'd775160064257445628},
        {64'd1098924405216917470},
        {64'd1863781237603223624},
        {64'd790381729229766398},
        {64'd1098924405216917470},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd1114415427349275283},
        {64'd808847097277379818},
        {64'd596828589218337826},
        {64'd330760979614274049},
        {64'd4349803816458794555},
        {64'd578739077902242850},
        {64'd330760979614274049},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd756201162802962713},
        {64'd66690625433381491},
        {64'd611682246103484322},
        {64'd1149941352894657557},
        {64'd1022963664536488677},
        {64'd544991620670102831},
        {64'd1149941352894657557},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd773999298348622632},
        {64'd441919094460623031},
        {64'd1036431620476294871},
        {64'd265266940119002720},
        {64'd2541675676191114756},
        {64'd441919094460623031},
        {64'd265266940119002720},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd632352089659195441},
        {64'd554433922346467269},
        {64'd651289513088373809},
        {64'd327484678248070126},
        {64'd2850087779045064517},
        {64'd72506280689865729},
        {64'd327484678248070126},
        {1'd0}
      },
      {
        {1'd0},
        {4'd6},
        {64'd751316387975571384},
        {64'd617128871946462362},
        {64'd788216112006338030},
        {64'd1094167526899186676},
        {64'd3219831875761420832},
        {64'd18140792658816702970},
        {64'd1094167526899186676},
        {1'd0}
      },
      {
        {1'd1},
        {4'd2},
        {64'd341603046690385513},
        {64'd23308969483731041},
        {64'd482255511267226920},
        {64'd506284367082604715},
        {64'd434838924625309677},
        {64'd505564480750957961},
        {64'd506284367082604715},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd1126722819440425677},
        {64'd817278496387404262},
        {64'd859555999965542145},
        {64'd1050246230107018792},
        {64'd4395836804990042725},
        {64'd812196183182151936},
        {64'd1050246230107018792},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd769930540971366242},
        {64'd64524193227225564},
        {64'd1072095771642353551},
        {64'd501957815896512795},
        {64'd1028027313880268498},
        {64'd495476670316155147},
        {64'd501957815896512795},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd773588673680130839},
        {64'd577925339242301887},
        {64'd206715480886209},
        {64'd244397469548096154},
        {64'd3085290030649338387},
        {64'd244599786440747995},
        {64'd244397469548096154},
        {1'd0}
      },
      {
        {1'd0},
        {4'd2},
        {64'd931422305862138371},
        {64'd118104809773309303},
        {64'd480201254464423231},
        {64'd255582357342028288},
        {64'd1403841544955375583},
        {64'd735783611806451519},
        {64'd255582357342028288},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd795151317050427103},
        {64'd896594382850788258},
        {64'd859709892774827999},
        {64'd257954227047318793},
        {64'd4381528848453580135},
        {64'd257954227047318793},
        {64'd257954227047318793},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd175959455021676869},
        {64'd361013055948620380},
        {64'd680350140418789899},
        {64'd455743996413491195},
        {64'd1620011678816158389},
        {64'd319337084470169519},
        {64'd455743996413491195},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd90481000911880086},
        {64'd501399981804029441},
        {64'd830666978375767898},
        {64'd1148982167232943188},
        {64'd2096080928127997850},
        {64'd1150422554116986718},
        {64'd1148982167232943188},
        {1'd0}
      },
      {
        {1'd1},
        {4'd7},
        {64'd502455366257286809},
        {64'd960623565581571380},
        {64'd150766284046204269},
        {64'd245757065567670743},
        {64'd4344949628583572329},
        {64'd960623565581571380},
        {64'd245757065567670743},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd930113865311746369},
        {64'd175070890352369345},
        {64'd514366262230445379},
        {64'd805759489908924528},
        {64'd1630397426721223749},
        {64'd1094346121796119923},
        {64'd805759489908924528},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd57884158320833968},
        {64'd33012865495543962},
        {64'd584371396828855280},
        {64'd849157567541524696},
        {64'd189935620303009816},
        {64'd5638296447299728},
        {64'd849157567541524696},
        {1'd0}
      },
      {
        {1'd1},
        {4'd6},
        {64'd231763707496170526},
        {64'd194636213789072862},
        {64'd129044885380461830},
        {64'd388533391995974300},
        {64'd1010308562652461974},
        {64'd18381152745300940584},
        {64'd388533391995974300},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd498530363177195850},
        {64'd474071177116854641},
        {64'd1016341751447247236},
        {64'd138864450208880668},
        {64'd2394815071644614414},
        {64'd138864450208880668},
        {64'd138864450208880668},
        {1'd0}
      },
      {
        {1'd1},
        {4'd0},
        {64'd519002793971381092},
        {64'd669506337717446578},
        {64'd653892412109155505},
        {64'd355273758432405838},
        {64'd3197028144841167404},
        {64'd649099055984829616},
        {64'd355273758432405838},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd698487305873808864},
        {64'd311958698635094234},
        {64'd115078982461317651},
        {64'd237940250836394761},
        {64'd1946322100414185800},
        {64'd74402996231365121},
        {64'd237940250836394761},
        {1'd0}
      },
      {
        {1'd0},
        {4'd1},
        {64'd465193278867515831},
        {64'd320532022240255113},
        {64'd388806280189807710},
        {64'd690940230277323271},
        {64'd1747321367828536283},
        {64'd1006545149321797215},
        {64'd690940230277323271},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd22399568880255913},
        {64'd267028626444729741},
        {64'd13289495247481252},
        {64'd543423807757741301},
        {64'd1090514074659174877},
        {64'd2850005733894308},
        {64'd543423807757741301},
        {1'd0}
      },
      {
        {1'd0},
        {4'd0},
        {64'd244252727490605211},
        {64'd1010685959893837610},
        {64'd364363167225850888},
        {64'd1152699804220354030},
        {64'd4286996567065955651},
        {64'd364283991038307336},
        {64'd1152699804220354030},
        {1'd0}
      },
      {
        {1'd0},
        {4'd7},
        {64'd110971566495168199},
        {64'd555425477363541999},
        {64'd169698942068938542},
        {64'd199292524206157032},
        {64'd2332673475949336195},
        {64'd199292524206157032},
        {64'd199292524206157032},
        {1'd0}
      }
    };

    // First reset test bench creation
    reset_tb = 1;
    #27ns reset_tb = 0;
  end

  always @(negedge clk) begin
    // Check test executed on positive edge of clk
    if (~reset_tb) begin
      if({PCBranch_E, aluResult_E, writeData_E, zero_E} !== {PCBranch_E_expected, aluResult_E_expected, writeData_E_expected, zero_E_expected}) begin
        $display("Error in test number %d with \
            input = { AluSrc = %d, AluControl = %b, PC_E = %d, signImm_E = %d, readData1_E = %d, readData2_E = %d } and \
            output = { PCBranch_E = %d, aluResult_E = %d, writeData_E = %d, zero_E = %d } --> \
            The expected output was { PCBranch_E_expected = %d, aluResult_E_expected = %d, writeData_E_expected = %d, zero_E_expected = %d }\
            ", test_number, AluSrc, AluControl, PC_E, signImm_E,
                 readData1_E, readData2_E, PCBranch_E, aluResult_E, writeData_E, zero_E,
                 PCBranch_E_expected, aluResult_E_expected, writeData_E_expected, zero_E_expected);
        cnt_errors++;
      end
      test_number++;

      if (test_number === CNT_TESTS) begin
        $display("%d tests completed with %d errors", CNT_TESTS, cnt_errors);
        #5ns $stop;
      end
    end

    // Prepare next test to positive edge of clk
    #2ns;
    {AluSrc, AluControl, PC_E, signImm_E, readData1_E, readData2_E, PCBranch_E_expected, aluResult_E_expected, writeData_E_expected, zero_E_expected} = test[test_number];
    #2ns;
  end

endmodule
